library verilog;
use verilog.vl_types.all;
entity main_tb is
end main_tb;
